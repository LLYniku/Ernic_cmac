


localparam [64*142-1 :0] reg_config = {
{32'h50060840, 32'h004c0387}, //142
{32'h50060844, 32'h04ffffb5},
{32'h50060884, 32'h008f503b},
{32'h50060804, 32'hcea61326}, //139
{32'h50060810, 32'h00608000},
{32'h5006083c, 32'h00400100},
{32'h50060848, 32'h00000007},
{32'h50060818, 32'h00140800},
{32'h50060888, 32'h70004f00}, //134
{32'h50060820, 32'h0fff001c},
{32'h50060800, 32'h045c0407},
{32'h50060828, 32'h0fff101c},
{32'h50060808, 32'h02040000},
{32'h50060850, 32'he2f8a222}, //129
{32'h50060854, 32'h0000e2de},
{32'h50060860, 32'h7481e444},
{32'h5006086c, 32'h3e52e18c},
{32'h50060864, 32'h780e5bcb},
{32'h50060868, 32'h5a95ddd8}, //124
{32'h50060740, 32'h00f9a408},
{32'h50060744, 32'h04ffff84},
{32'h50060784, 32'h007f503b},
{32'h50060704, 32'h167b4025},
{32'h50060710, 32'h00607000}, //119
{32'h5006073c, 32'h00800040},
{32'h50060748, 32'h00000006},
{32'h50060718, 32'h00140700},
{32'h50060788, 32'h70003f00},
{32'h50060720, 32'h0fff0018}, //114
{32'h50060700, 32'h012b0427},
{32'h50060728, 32'h0fff1018},
{32'h50060708, 32'h02038000},
{32'h50060750, 32'had424e4e},
{32'h50060754, 32'h000002dd}, //109
{32'h50060760, 32'h4abea0cf},
{32'h5006076c, 32'h00897117},
{32'h50060764, 32'h6bb328b7},
{32'h50060768, 32'hd52a10d0},
{32'h50060640, 32'h0000000a}, //104
{32'h50060644, 32'h04000001},
{32'h50060684, 32'h006f503b},
{32'h50060604, 32'h50e92b2a},
{32'h50060610, 32'h00606000},
{32'h5006063c, 32'h00400040},  //99
{32'h50060648, 32'h00000005},
{32'h50060618, 32'h00140600},
{32'h50060688, 32'h70002f00},
{32'h50060620, 32'h0fff0014},
{32'h50060600, 32'h02940407},  //94
{32'h50060628, 32'h0fff1014},  
{32'h50060608, 32'h02030000},  
{32'h50060650, 32'h27fbffe6},  
{32'h50060654, 32'h00008b09},  
{32'h50060660, 32'h98b129af},  //89
{32'h5006066c, 32'h8aa47e41},  
{32'h50060664, 32'h2ee66645},  
{32'h50060668, 32'h02c1bf38},  
{32'h50060540, 32'h00974470},  
{32'h50060544, 32'h04c02aa9},  //84
{32'h50060584, 32'h005f503b},  
{32'h50060504, 32'h9ff2b002},  
{32'h50060510, 32'h00800000},  
{32'h5006053c, 32'h00500200},  
{32'h50060548, 32'h00000004},  //79
{32'h50060518, 32'h00360000},  
{32'h50060588, 32'h70001f00},  
{32'h50060520, 32'h1ffff010},  
{32'h50060500, 32'h06f80407},  
{32'h50060528, 32'h2fff1010},   //74
{32'h50060508, 32'h04000000},  
{32'h50060550, 32'h60660f2e},  
{32'h50060554, 32'h000016e4},  
{32'h50060560, 32'h622c6007},  
{32'h5006056c, 32'hcebceaf4},   //69
{32'h50060554, 32'h9840f9eb},  
{32'h50060568, 32'h460a5e88},  
{32'h50060340, 32'h00774470},  
{32'h50060344, 32'h04a02aa9},  
{32'h500600a0, 32'h0c000000},   //64
//{32'h50060030, 32'h00100000},  //UNKNOWN 1
{32'h50060010, 32'h00112233},  //63
{32'h50060070, 32'hc0a8010c},  //62 IPv4 address 
{32'h50060014, 32'h00004455},  //61
{32'h50060024, 32'hac92135d},  //60
{32'h50060028, 32'h013248eb},  //59
{32'h500600a8, 32'h10000080},  //58
{32'h50060020, 32'hf38590ba},  //57// IPv6 address
{32'h5006002c, 32'hafb1f367},  //56
//{32'h50060038, 32'h00800080},  //UNKNOWN 2
{32'h50060068, 32'h01000040},  //55
//{32'h50060048, 32'h00400100},  //UNKNOWN 4
//{32'h50060058, 32'h02000020},    //UNKNOWN 6
{32'h50060060, 32'h00110000},  //54
//{32'h50060050, 32'h00120000},  //UNKNOWN 5
//{32'h50060040, 32'hb4000000},  //UNKNOWN 3
{32'h50060210, 32'h0b000000},  //53
{32'h5006023c, 32'h00800040},  //52
{32'h50060248, 32'h00000001},  //51
{32'h50060218, 32'h0b800000},  //50
{32'h50060220, 32'h0fff0000},  //49
{32'h50060200, 32'h024f0435},  //48
{32'h50060250, 32'hd1677ed7},  //47
{32'h50060254, 32'h0000c918},  //46
{32'h50060228, 32'h0fff1000},  //45
{32'h50060208, 32'h08000000},  //44
{32'h50060260, 32'ha3c9ba8b},  //43
{32'h5006026c, 32'h6f2a46fe},  //42
{32'h50060264, 32'h823b88db},  //41 
{32'h50060268, 32'h1798f443},  //40
{32'h50060384, 32'h004e503b},  //39
{32'h50060304, 32'h9bf1b002},  //38
{32'h50060310, 32'h00600000},  //37
{32'h5006033c, 32'h00400100},  //36
{32'h50060348, 32'h00000002},  //35
{32'h50060318, 32'h00140000},  //34
{32'h50060388, 32'h70000600},  //33
{32'h50060320, 32'h0fff0004},  //32
{32'h50060300, 32'h04f80407},  //31
{32'h50060328, 32'h0fff1004},  //30
{32'h50060308, 32'h02000000},  //29
{32'h50060484, 32'h00d47c2d},  //28
{32'h50060488, 32'h70000600},  //27
{32'h50060440, 32'h00e21df7},  //26
{32'h50060444, 32'h040b77ce},  //25
{32'h50060350, 32'h50560f2e},  //24
{32'h50060354, 32'h000016c4},  //23
{32'h50060360, 32'h610c6007},  //22
{32'h5006036c, 32'hccbceaf4},  //21
{32'h50060364, 32'h9640f9eb},  //20
{32'h50060368, 32'h440a5e88},  //19
{32'h50060404, 32'hd836ba10},  //18
{32'h50060410, 32'h00604000},  //17
{32'h5006043c, 32'h00400100},  //16
{32'h50060448, 32'h00000003},  //15
{32'h50060418, 32'h00140400},  //14
{32'h50060420, 32'h0fff0008},  //13
{32'h50060400, 32'h01dd030b},  //12
{32'h50060428, 32'h0fff1008},  //11
{32'h50060408, 32'h02010000},  //10
{32'h50060000, 32'he3480789},  //9
{32'h50060180, 32'h00000070},  //8
{32'h50060450, 32'hddf1c650},  //7
{32'h50060454, 32'h00006b4b},  //6
{32'h50060460, 32'hc0a81621},  //5
{32'h5006046c, 32'he9a855a0},  //4
{32'h50060464, 32'h92e8a89f},  //3
{32'h50060468, 32'h28640e94},  //2
{32'h50060000, 32'he348078b}}; //1




localparam [16*512-1:0] rdma_rdwr_wqe = {
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6161c8ce364edf276000e6a8010000000100000000008c00F0000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6161c7ce364edf276000e6a8010000000100000000008c00E0000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6161c6ce364edf276000e6a8010000000100000000008c00D0000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6161c5ce364edf276000e6a8010000000100000000008c00C0000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6161c4ce364edf276000e6a8010000000100000000008c00B0000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6161c3ce364edf276000e6a8010000000100000000008c00A0000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6161c2ce364edf276000e6a8010000000100000000008c0090000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6161c1ce364edf276000e6a8010000000100000000008c0080000000e0a6},// RDMA wr wqe starts
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6140a5ce364edf276000e6a8010400000100000000008c0070000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6140a5ce364edf276000e6a8010400000100000000008c0060000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6140a5ce364edf276000e6a8010400000100000000008c0050000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6140a5ce364edf276000e6a8010400000100000000008c0040000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6140a5ce364edf276000e6a8010400000100000000008c0030000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6140a5ce364edf276000e6a8010400000100000000008c0020000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6140a5ce364edf276000e6a8010400000100000000008c0010000000e0a6},
{512'h0000000000000000000000000000000000000000000000000000000000000000d30e6140a5ce364edf276000e6a8010400000100000000008c0000000000e0a6} // RDMA rd wqe starts
};

localparam NUM_RD_WQE = 8;
localparam NUM_WR_WQE = 8;

localparam EN_SEND_PKT = 1;
localparam EN_RDMA_WR_PKT =  1;
localparam EN_RDMA_RD_PKT = 1;


//target code ends
//initiator code

